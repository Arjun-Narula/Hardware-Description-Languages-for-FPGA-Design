LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ALU IS
PORT( Op_code : IN STD_LOGIC_VECTOR( 2 DOWNTO 0 );
A, B : IN STD_LOGIC_VECTOR( 31 DOWNTO 0 );
Y : OUT STD_LOGIC_VECTOR( 31 DOWNTO 0 ) );
END ALU;
ARCHITECTURE ARCH_ALU OF ALU IS
BEGIN
Y<=A WHEN (OP_CODE = "000") ELSE
   A+B WHEN (OP_CODE = "001") ELSE
   A-B WHEN (OP_CODE = "010") ELSE
   A AND B WHEN (OP_CODE = "011") ELSE
   A OR B WHEN (OP_CODE = "100") ELSE
   A+1 WHEN (OP_CODE = "101") ELSE
   A-1 WHEN (OP_CODE = "110") ELSE
   B WHEN (OP_CODE = "111") ELSE
   "00000000000000000000000000000000";
END ARCH_ALU;
